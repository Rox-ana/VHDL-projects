-------------------------------------------------------------------------------
--
-- Title       : ROM
-- Design      : coDesignCPU
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : ROM.vhd
-- Generated   : Sat Jun 16 19:46:57 2018
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {ROM} architecture {ROM}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
entity ROM is
	port(
	mem_out : out std_logic_vector(5 downto 0);
	RD : in std_logic; 
	
	mem_in : in std_logic_vector(5 downto 0)
	);
end ROM;

--}} End of automatically maintained section

architecture ROM of ROM is

type memory is array(63 downto 0) of std_logic_vector(5 downto 0);
constant mem : memory := (
0 => "000000",
1 => "000101",
2 => "000100",
3 => "000110",
4 => "001000",
5 => "000000",
6 => "001100",
7 => "000001",
8 => "011000",
9 => "100111",
10 => "110100",
11 => "001000",
12 => "000000",
13 => "000111",
14 => "000100",
15 => "001000",
16 => "001000",
17 => "000000",
18 => "001100",
19 => "000000",
20 => "011000",
21 => "011101",
22 => "010001",
23 => "010110",
24 => "100010",
25 => "100111",
26 => "000000",
27 => "000101",
28 => "000100",
29 => "001001",
30 => "100100",
31 => "001000",
32 => "000001",
33 => "001100",
34 => "000000",
35 => "011100",
36 => "100110",
37 => "010011",
38 => "110100",
39 => "100100",
40 => "000000",
41 => "001111",
42 => "000100",
43 => "010100",
44 => "001000",
45 => "000000",
46 => "011000",
47 => "010001",
48 => "100110",
49 => "000000",
50 => "000000",
51 => "000000",
52 => "000000",
53 => "000000",
54 => "000000",
55 => "000000",
56 => "000000",
57 => "000000",
58 => "000000",
59 => "000000",
60 => "000000",
61 => "000000",
62 => "000000",
63 => "000000"
);

begin
	
	 mem_out <= Mem(to_integer(unsigned(mem_in))) when rd = '1' else (others => 'Z'); 
	

end ROM;
